package dma_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "dma_sequence_item.sv"  
  //REGISTER CONFIGURATION FILES
  `include "registers/config_reg.sv"
  `include "registers/ctrl_reg.sv" 
  `include "registers/descriptor_addr_reg.sv"
  `include "registers/error_status_reg.sv"
  `include "registers/extra_info_reg.sv"
  `include "registers/intr_reg.sv"
  `include "registers/io_addr_reg.sv"
  `include "registers/mem_addr_reg.sv"
  `include "registers/status_reg.sv"
  `include "registers/transfer_count_reg.sv"

  `include "dma_reg_block.sv"
  `include "dma_adapter.sv"        

  //ALL SEQUENCES
  `include "tests/sequences/dma_sequence.sv"
  `include "tests/sequences/reset_all_sequence.sv"
  `include "tests/sequences/config_sequence.sv"
  `include "tests/sequences/ctrl_sequence.sv"
  `include "tests/sequences/descriptor_addr_sequence.sv"
  `include "tests/sequences/error_status_sequence.sv"
  `include "tests/sequences/extra_info_sequence.sv"
  `include "tests/sequences/intr_sequence.sv"
  `include "tests/sequences/io_addr_sequence.sv"
  `include "tests/sequences/mem_addr_sequence.sv"
  `include "tests/sequences/status_sequence.sv"
  `include "tests/sequences/transfer_count_sequence.sv"
  `include "tests/sequences/regression_sequence.sv"

  `include "dma_monitor.sv"        
  `include "dma_driver.sv"         
  `include "dma_sequencer.sv"
  `include "dma_agent.sv"           
  `include "dma_subscriber.sv"
  `include "dma_environment.sv"   
  `include "dma_report_server.sv"   

  //ALL TESTS
  `include "tests/config_test.sv"
  `include "tests/ctrl_test.sv"
  `include "tests/descriptor_addr_test.sv"
  `include "tests/error_status_test.sv"
  `include "tests/extra_info_test.sv"
  `include "tests/intr_test.sv"
  `include "tests/io_addr_test.sv"
  `include "tests/mem_addr_test.sv"
  `include "tests/reset_all_test.sv"
  `include "tests/status_test.sv"
  `include "tests/transfer_count_test.sv"
  `include "tests/regression_test.sv"
endpackage
