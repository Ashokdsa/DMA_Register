`include "uvm_macros.svh"
import uvm_pkg::*;

package dma_reg_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
//  `include "dma_register.sv"
endpackage
